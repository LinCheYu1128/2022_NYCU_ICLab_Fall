//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//      (C) Copyright NCTU OASIS Lab      
//            All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2022 ICLAB fall Course
//   Lab05			: SRAM, Matrix Multiplication with Systolic Array
//   Author         : Jia Fu-Tsao (jiafutsao.ee10g@nctu.edu.tw)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : TESTBED.v
//   Module Name : TESTBED
//   Release version : v1.0
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################
`ifdef RTL
	`timescale 1ns/10ps
	`include "MMSA.v"
	`define CYCLE_TIME 20.0
`endif
`ifdef GATE
	`timescale 1ns/10ps
	`include "MMSA_SYN.v"
	`define CYCLE_TIME 20.0
`endif

module PATTERN(
// output signals
    clk,
    rst_n,
    in_valid,
	in_valid2,
    matrix,
    matrix_size,
    i_mat_idx, 
    w_mat_idx,
// input signals
    out_valid,
    out_value
);
//================================================================
//   INPUT AND OUTPUT DECLARATION                         
//================================================================
output reg 		  clk, rst_n, in_valid, in_valid2;
output reg [15:0] matrix;
output reg [1:0]  matrix_size;
output reg [3:0]  i_mat_idx, w_mat_idx;

input 				out_valid;
input signed [39:0] out_value;
//================================================================
//   parameters & integers
//================================================================
integer ans_count, cycles, total_cycles;
integer patcount, PATNUM;
integer in_read, out_read;
integer i, j, k, a, gap;

integer temp_cycle;
integer img_size, matrix_num, out_size;
integer idx_x[0:15];
integer idx_w[0:15];
//================================================================
//    wires % registers
//================================================================
reg signed [39:0] y_temp[0:30];
//================================================================
//    clock
//================================================================
always	#(`CYCLE_TIME/2.0) clk = ~clk;
initial	clk = 0;
//================================================================
//    initial
//================================================================
initial begin
    in_read = $fopen("../00_TESTBED/input.txt", "r");
	out_read = $fopen("../00_TESTBED/output.txt", "r");
	a = $fscanf(in_read, "%d\n", PATNUM);

    rst_n       = 1'b1;
    in_valid    = 1'b0;
	in_valid2   = 1'b0;
    matrix      = 16'bx;
    matrix_size = 2'bx;
    i_mat_idx   = 4'bx;
    w_mat_idx   = 4'bx;

    total_cycles = 0;
	reset_task;

    for(patcount = 0; patcount < PATNUM; patcount = patcount+1)begin
		input_matrix_task;
        a = $fscanf(out_read, "%d\n", out_size);
        temp_cycle = 0;
        for(matrix_num=0; matrix_num<16; matrix_num=matrix_num+1)begin  
            input_idx_task;
            wait_outvalid_task;
            check_ans_task;
        end
		$display("\033[0;34mPASS PATTERN NO.%4d,\033[m \033[0;32mexecution cycle : %3d\033[m",patcount ,temp_cycle);
	end
	YOU_PASS_task;
end

task check_ans_task ; begin
    ans_count = 0;
    for(i=0; i < out_size; i=i+1)begin
		a = $fscanf(out_read, "%d\n", y_temp[i]);
	end
    while (out_valid === 1) begin
        if(ans_count >= out_size)begin
			$display ("----------------------------------------------------------------------------------------------------------------------");
			$display ("                                             The out_valid should be %d cycles                               ",out_size);
			$display ("----------------------------------------------------------------------------------------------------------------------");
			$finish;
		end
        else begin
            if(y_temp[ans_count] !== out_value )begin
                $display ("----------------------------------------------------------------------------------------------------------------------");
				$display ("                                                  Your Answer is Wrong!             						             ");
				$display ("                                                  Your Answer is : %d       	                               ",out_value);
				$display ("                                               Correct Answer is : %d          			           ",y_temp[ans_count]);
				$display ("----------------------------------------------------------------------------------------------------------------------");
				$finish;
            end
            ans_count = ans_count+1;
        end
        @(negedge clk);
    end
    if(ans_count!=out_size)begin
		$display ("----------------------------------------------------------------------------------------------------------------------");
        $display ("                                             The out_valid should be %d cycles                               ",out_size);
        $display ("----------------------------------------------------------------------------------------------------------------------");
        $finish;
	end
end endtask

task input_idx_task ; begin
    i_mat_idx = idx_x[matrix_num];
    w_mat_idx = idx_w[matrix_num];
    in_valid2 = 1'b1;
    @(negedge clk);
    i_mat_idx = 'bx;
    w_mat_idx = 'bx;
    in_valid2 = 1'b0;
end endtask

task input_matrix_task ; begin
    gap = $urandom_range(1,5);
	repeat(gap) @(negedge clk);
    a = $fscanf(in_read, "%d\n", img_size);
    
    for(i=0; i<32; i=i+1)begin
        for(j=0; j<img_size; j=j+1)begin
            for(k=0; k<img_size; k=k+1)begin
                if(i==0 && j==0 && k==0)begin
                    if(img_size==2) matrix_size = 2'b00;
                    else if(img_size==4) matrix_size = 2'b01;
                    else if(img_size==8) matrix_size = 2'b10;
                    else matrix_size = 2'b11;
                end
                else matrix_size = 2'bx;
                in_valid = 1'b1;
                a = $fscanf(in_read, "%d\n", matrix);
                @(negedge clk);
            end
        end
    end
    matrix      = 16'bx;
    in_valid    = 1'b0;
    @(negedge clk);
    for(i=0; i<16; i=i+1)begin
        a = $fscanf(in_read, "%d\n", idx_x[i]);
    end
    for(i=0; i<16; i=i+1)begin
        a = $fscanf(in_read, "%d\n", idx_w[i]);
    end
end endtask

task wait_outvalid_task ; begin
	cycles = 0 ;
	while( out_valid === 0 ) begin
		cycles = cycles + 1 ;
        temp_cycle = temp_cycle + 1;
		if (cycles==2000) begin 
			$display ("----------------------------------------------------------------------------------------------------------------------");
			$display ("                                             Exceed maximun cycle!!!                                                  ");
			$display ("----------------------------------------------------------------------------------------------------------------------");
			$finish;
		end
		@(negedge clk);
	end
	total_cycles = total_cycles + cycles ;
end endtask

task reset_task ;  begin
	force clk = 0;
	#(20); rst_n = 0;
	#(20);
	if((out_valid!==0) || (out_value!==0))begin
		reset_fail;
	end
	#(20);rst_n = 1;
	#(6); release clk;
end endtask

always @(negedge clk) begin
  if(out_valid === 0 && out_value !== 0)begin
    $display ("----------------------------------------------------------------------------------------------------------------------");
	$display ("                                          out should be 0 when out_valid is low         						         ");
	$display ("----------------------------------------------------------------------------------------------------------------------");
	$finish;
  end
end

always @(negedge clk) begin
  if((in_valid === 1 || in_valid2 === 1) && out_valid !== 0)begin
    $display ("----------------------------------------------------------------------------------------------------------------------");
	$display ("                                     out_valid should not be high when in_valid is high 						         ");
	$display ("----------------------------------------------------------------------------------------------------------------------");
	$finish;
  end
end

task reset_fail ; begin
	$display ("----------------------------------------------------------------------------------------------------------------------");
	$display ("                                                  Oops! Reset is Wrong                						         ");
	$display ("----------------------------------------------------------------------------------------------------------------------");
	$finish;
end endtask

task YOU_PASS_task; begin                                                                                                                                                                                            
    $display("\033[1;32m                                          .:---:.                                                                         ");                                  
    $display("\033[1;32m                                       .*aa&&&&&aa#=                                                                      ");                                  
    $display("\033[1;32m                                    .#a#*+***###&aaaa&&&&&##**+=-::.                                                      ");                                  
    $display("\033[1;32m                                 .=*&aa&####***++++++++++++++****##&&&&##+=-:                                             ");                                  
    $display("\033[1;32m                              :*&aa&#*+++++++++++++++++++++++++++++++++++*##&&&#+=:.                                      ");                                  
    $display("\033[1;32m                           :+aa&*+=====================+++++++++++++++++++++++++*##&&#+-.                                 ");                                  
    $display("\033[1;32m                         =&a#*================================+++++++++++++++++++++++*#&a&*=.                             ");                                  
    $display("\033[1;32m                       +aa*===============+&&+==================++==+++++++++++++++++++++*#&aa*-     .----.               ");                                  
    $display("\033[1;32m                     =a&*==================**==================+aa+=====+++++++++++++++++++++#&aa#=+aa####&&&*-           ");                                  
    $display("\033[1;32m                   .&a*======================================================+++++++++++++++++++*&aa*++++++++*&a*.        ");                                  
    $display("\033[1;32m                  :a&+===========================================================++++++++++++++++++*++++*###**++#a*       ");                                  
    $display("\033[1;32m                 :a&==============++**#######*#aa*****#####**++=====================+++++++++++++++++++&a&&&&a&#++&&.     ");                                  
    $display("\033[1;32m                 &a=========+*#&#*+-:.       \033[1;37m=*::#:        .:-=#a&##*+\033[1;32m=================+++++++++++++++*a&&&&&&&a&++&&");                                  
    $display("\033[1;32m                =a+=====+*#*=:\033[1;37m***=         -*-   \033[1;37m.*+         =*=.:#:.\033[1;32m-=+*#*+==============+++++++++++++&&&&&&&&&&+++a*");                                  
    $display("\033[1;32m                #a===*##=.   \033[1;37m-##  #+     :*= \033[1;32m::    \033[1;37m=#.    .+*:    \033[1;32m.\033[1;37m#:     \033[1;32m.-+*#*+============+++++++++++#&a&&&a&*+++&a");                                  
    $display("\033[1;32m                #a*&*+#*\033[1;37m=   .&. \033[1;32m#+:\033[1;37m:*+.-*=  \033[1;32m*&*    \033[1;37m :*= -*+.     \033[1;32m.:.\033[1;37m#-         \033[1;32m.=+#*+===========+++++++++++*#**+++++&&");                                  
    $display("\033[1;32m                =a&. #- \033[1;37m-*-:#.\033[1;32m.#+-*  \033[1;37m.=: \033[1;32m .#-+*      \033[1;37m -+-        \033[1;32m-a. \033[1;37m*+        \033[1;32m:++=:a*#*+=========+++++++++++++++++#a-");                                  
    $display("\033[1;32m                 &a::#   \033[1;37m -=. \033[1;32m*+*&+      .#: =*..               :+a=  \033[1;37m=*    -++-.-  -* \033[1;32m:=*#+========+++++++++++++#a#.");                                  
    $display("\033[1;32m                 :aa#:       *&#:&:      *=  :&&#...           ::##+   \033[1;37m:*+++:        *=   \033[1;32m:=*#+========+++++++++++&a:  ");                                  
    $display("\033[1;32m                .#&:.       =a- .a-+*##**#*-  #*=#+++==--:::::::-a-*     .-=---+*=*  \033[1;37m#&:     \033[1;32m.=#*========++++++++++&&  ");                                  
    $display("\033[1;32m               =a#.        :&. :*a*-. .           ..::--=++++++*#+-*     .--=+&&#&&:++\033[1;37m.&.      \033[1;32m.*a*========++++++++*a+ ");                                  
    $display("\033[1;32m             -&&- :*      .&:.##-:=*******=.                      .=+++++++++*+  .-*a+.\033[1;37m:#:-=*++-:+*\033[1;32m#*=======++++++++&a ");                                  
    $display("\033[1;32m            #a&===&:      ++ &-.*#-:.....:+&-                            .-*##**+=:  =&+.-:.&    \033[1;37m:& \033[1;32m-#+=======++++++*a-");                                  
    $display("\033[1;32m             .:-#a+      .&.   &+..........:&-                         :*#+-:...:-+&-  +*   a.    \033[1;37m#- \033[1;32m &+=======++++++a+");                                  
    $display("\033[1;32m                a&.      ++   -&          ..&=                        :a+..........:a:      a.    \033[1;37m:#  \033[1;32m:&========+++++a*");                                  
    $display("\033[1;32m               =a-      .&.   -&           +#.              .         =&         ...*+      a:     \033[1;37m#: \033[1;32m.&*========++++a*");                                  
    $display("\033[1;32m               &&       =#     +#:      :+&=       +:==.  -##*        :a.           &-      a:     \033[1;37m:+=-\033[1;32m+#=========+++a*");                                  
    $display("\033[1;32m              .a+      .#-   \033[1;31m...-+#****#*=.        \033[1;32m.+#=#+**--&         -&+:       -#+      :&:.        :a=========++*a=");                                  
    $display("\033[1;32m              =a:     .:a. \033[1;31m......:..........        \033[1;32m-*:------&       \033[1;31m....-*#******+:     \033[1;32m##+*:.  .=:   .a==========+#a:");                                  
    $display("\033[1;32m              *a.     :-&  \033[1;31m....:=:...:-:.....       \033[1;32m=*-------&      \033[1;31m......::.....:...   \033[1;32m-#:#*-:=*+*+    a==========+&& ");                                  
    $display("\033[1;32m           --:*&     .:+*  \033[1;31m...:=:...:=:......       \033[1;32m=*------+*      \033[1;31m.....--:...:-:.... \033[1;32m.#&#####&*=+=   .a==========+a= ");                                  
    $display("\033[1;32m          .a&aa&     ::*=   \033[1;31m...:....::......        \033[1;32m-*------#=      \033[1;31m....::....--......\033[1;32m+&*+++++==+#a:   :&==========&&  ");                                  
    $display("\033[1;32m           a*=&a+-.  ::*=..   \033[1;31m....:........         \033[1;32m:#:-----a.       \033[1;31m................\033[1;32m##++++=======&-   =#=========+a-  ");                                  
    $display("\033[1;32m           aa*+++*##-::*&*::    \033[1;37m.:++:.           .   \033[1;32m&-----+*           \033[1;31m.:-=::....  \033[1;32m+#+++=========**   **=========a*   ");                                  
    $display("\033[1;32m       .=*aa+====+++##\033[1;37m+#:-#:: .:=#.:#+:.      .:+*-..\033[1;32m=*----&- \033[1;37m+++-:.     :+*-+*=..  \033[1;32m.a+++==========**   &+========#a.  ");                                  
    $display("\033[1;32m      .aa--a=======++\033[1;37m*&.  *+:::#=    =#-:.   .-#- =*=.\033[1;32m+*=+#+\033[1;37m-# .=*+-:. :=#    -**:\033[1;32m.#*++===========**  :&========#a:    ");                                  
    $display("\033[1;32m       .#a+a========*\033[1;37m&.    &-=#:      .*+:..:=#.    -#=:\033[1;32m---\033[1;37m&:     .+*=:-&       .+\033[1;32m#&++============#-  **=======#a-     ");                                  
    $display("\033[1;32m         :#a*======+a#*+=-:\033[1;37m=&*          -#-:*+        -#=:&:         -*&-..:-\033[1;32m=++*#a*++===========+&--.a=======#a:");                                  
    $display("\033[1;32m           +a+======#&*==++*#***++==-::..\033[1;37m:##=           +&=..\033[1;32m::--=+++**##**++====+&++============&+&.+#=====+&&. ");                                  
    $display("\033[1;32m            =a*=======#&*===========+++****#***********#*****++++================&*+============#*#+:&=====#a=     ");                                  
    $display("\033[1;32m             :&&+=======#&#+====================================================+&++===========*&&###+===*a*.      ");                                  
    $display("\033[1;32m              .aa#========*#&#+=================================================&*+===========+a&**a*==#a*.        ");                                  
    $display("\033[1;32m               &&*a#+=======+*#&#*+============================================*&+===========+a#+++\033[1;31m&#&aa-");                                  
    $display("\033[1;32m               -aa&*a&+=========+*#&##*+=======================================a+===========+&*+=\033[1;31m+a&&&&aa+");                                  
    $display("\033[1;32m                =+. +a*##+===========+***=====================================*#============&*+===\033[1;31ma&&&&&a-");                                  
    $display("\033[1;32m                     *a-#aa#*=+*=================---\033[1;33m:::::::::::::\033[1;32m---=======================*&+====\033[1;31m#a&&&aa#&&.            ");                                  
    $display("\033[1;32m                      *aa#.=#aa*============--\033[1;33m::::::::::::::::::::::::::\033[1;32m-==================++======\033[1;31m&&&aaa&&a*            ");                                  
    $display("\033[1;32m                       -*.   =a*=========-\033[1;33m::::::::::::::::::::::::::::::::::\033[1;32m-======================\033[1;31m+a&&&&&&a& .-+:       ");                                  
    $display("\033[1;32m                             -a+=======-\033[1;33m::::::::::::::::::::::::::::::::::::::\033[1;32m-=====================\033[1;31m+&&&&&&aa&aaaa:  :.  ");                                  
    $display("\033[1;32m                             .a#=====-\033[1;33m:::::::::::::::::::::::::::::::::::::::::::\033[1;32m=====================\033[1;31m#a&&&aa&&&&a&+&aa= ");                                  
    $display("\033[1;32m                              #&====\033[1;33m:::::::::::::::::::::::::::::::::::::::::::::::\033[1;32m-===================\033[1;31m+&&&&&&&&&aa&&&aa:");                                  
    $display("\033[1;32m                              :a*==\033[1;33m::::::::::::::::::::::::::::::::::::::::::::::::::\033[1;32m====================\033[1;31m+##&&&&&&&&&&##=");                                  
    $display("\033[1;34m      ===============================================================================================================");
	$display("\033[1;34m                                                  Congratulations!                						             ");
	$display("\033[1;34m                                           You have passed all patterns!          						             ");
	$display("\033[1;34m                                           Your execution cycles = %5d cycles   					   ", total_cycles);
	$display("\033[1;34m                                           Your clock period = %.1f ns        					        ", `CYCLE_TIME);
	$display("\033[1;34m                                           Your total latency = %.1f ns                    ", total_cycles*`CYCLE_TIME);
    $display("\033[1;34m      ===============================================================================================================");  
    $display("\033[1;0m"); 
    $finish;

end endtask

endmodule